//
//
//
 module Room_FSM (
	input clk, current, N, S, W, E,
	output next
 );

 
 endmodule
 